 module MIPS_SC(//);
 endmodule 